** Profile: "Esquematico-Realimentacion"  [ C:\Users\Emanuel\Desktop\DCE-Amplificador-Clase-D\Calculo de realimentador\PSpice\Amplificador Clase D-PSpiceFiles\Esquematico\Realimentacion.sim ] 

** Creating circuit file "Realimentacion.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "../../../libraries/phb27nq10t/phb27nq10t.lib" 
.LIB "../../../libraries/ucc20520_pspice_trans/ucc20520_trans.lib" 
* From [PSPICE NETLIST] section of C:\Users\Emanuel\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice\17.2.0\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 2m 0 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\Esquematico.net" 


.END
