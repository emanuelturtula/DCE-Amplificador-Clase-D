** Profile: "Esquematico-Transient"  [ C:\Users\Emanuel\Desktop\DCE-Amplificador-Clase-D\Amplificador\amplificador clase d-pspicefiles\esquematico\transient.sim ] 

** Creating circuit file "Transient.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "../../../libraries/phb27nq10t/phb27nq10t.lib" 
.LIB "../../../libraries/ucc20520_pspice_trans/ucc20520_trans.lib" 
* From [PSPICE NETLIST] section of C:\Users\Emanuel\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice\17.2.0\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 10ms 0 
.OPTIONS ADVCONV
.OPTIONS SPEED_LEVEL= 0
.AUTOCONVERGE ITL1=1000 ITL2=1000 ITL4=1000 RELTOL=0.05 ABSTOL=1.0E-6 VNTOL=.001 PIVTOL=1.0E-10 
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\Esquematico.net" 


.END
